localparam ABITS = 12;
localparam DBITS = 18;

localparam DEPTH = 2**ABITS;
